//List of Include Files

 `include "spi_base_test.sv"
 `include "reset_test.sv"
 `include "lsb_fst_data_test.sv"
 `include "msb_fst_data_test.sv"
 `include "miso_data_test.sv"


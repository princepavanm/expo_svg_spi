`include "reset_seq.sv"
`include "lsb_8bit_data.sv"
`include "lsb_16bit_data.sv"
`include "lsb_32bit_data.sv"
`include "lsb_64bit_data.sv"
`include "lsb_128bit_data.sv"
`include "msb_8bit_data_seq.sv"
`include "msb_16bit_data_seq.sv"
`include "msb_32bit_data_seq.sv"
`include "msb_64bit_data_seq.sv"
`include "msb_128bit_data_seq.sv"
`include "miso_data.sv"
`include "Rx_raising_Tx_falling_seq.sv"
`include "Rx_falling_Tx_raising_seq.sv"


`define CTRL_STATUS_ADDR     32'h 10
`define TX0_ADDR             32'h 00
`define RX0_ADDR             32'h 00
`define TX1_ADDR    	     32'h 04
`define RX1_ADDR    	     32'h 04
`define TX2_ADDR    	     32'h 08
`define RX2_ADDR    	     32'h 08
`define TX3_ADDR    	     32'h 0C
`define RX3_ADDR    	     32'h 0C
`define SS_ADDR              32'h 18
`define DIVIDER_ADDR         32'h 14


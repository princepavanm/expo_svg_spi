class wb_monitor extends uvm_monitor;

  `uvm_component_utils(wb_monitor)

  //virtual interface
  virtual wb_intf      wb_vif;

bit [63:0] packet;
bit [127:0] cntrl_status_reg;
  uvm_analysis_port #(wb_trans) wb_analysis_port;

  //wb transactor
  wb_trans   wb_trans_h;
 // int temp[5];
  /**********************constructor********************************/
  function new(string name, uvm_component parent);
    super.new(name,parent);
    wb_trans_h=new();
    wb_analysis_port = new("wb_analysis_port", this);
  endfunction 

/*********************build phase**********************/
 virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if (!uvm_config_db#(virtual wb_intf)::get(this,"*","wb_vif",wb_vif))
      `uvm_fatal("WB_DRV","**** Could not get virtual interface ****");
  endfunction: build_phase

/*******************run phase***********************/
virtual task run_phase(uvm_phase phase);
	
	wb_trans_h=wb_trans::type_id::create("wb_trans");
 	`uvm_info("WB_MON","WB Monitor Run Phase", UVM_LOW)

	`uvm_info("WB_MONITOR","WB_MONITOR_BEFORE_RAISE_OBJECTION ", UVM_HIGH)
	phase.raise_objection(this);
  	`uvm_info("WB_MONITOR","WB_MONITOR_AFTER_RAISE_OBJECTION ", UVM_HIGH)

	wait(wb_vif.rst==0);
	forever
	begin
     			@((wb_vif.clk) && !wb_vif.rst )
		 begin
		//	@(posedge wb_vif.clk);
		 //	if(wb_vif.wb_cyc_i == 1 && wb_vif.wb_stb_i == 1 && wb_vif.wb_sel_i == 111 && wb_vif.wb_ack_o==1) begin 
			wb_trans_h.wr_en <=  wb_vif.wb_we_i;

		if(wb_trans_h.wr_en==1)	begin	
			@(posedge wb_vif.clk);
			wb_trans_h.reg_addr    <= wb_vif.wb_adr_i;
			wb_trans_h.reg_wr_data <= wb_vif.wb_dat_i;

		
			if(wb_trans_h.reg_addr==`SS_ADDR) begin
				packet[31:0]=wb_trans_h.reg_wr_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h packet0=%h ",$time,wb_trans_h.reg_addr,packet[31:0]),UVM_HIGH)
			end

			if(wb_trans_h.reg_addr==`DIVIDER_ADDR) begin
				packet[63:32]=wb_trans_h.reg_wr_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h packet1=%h ",$time,wb_trans_h.reg_addr,packet[63:32]),UVM_HIGH)
			end

			if(wb_trans_h.reg_addr==`TX0_ADDR) begin
				wb_trans_h.mon_data[31:0]=wb_trans_h.reg_wr_data;
		//	`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_data0=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_data[31:0]),UVM_MEDIUM)
			end

			else if(wb_trans_h.reg_addr==`TX1_ADDR) begin
				wb_trans_h.mon_data[63:32]=wb_trans_h.reg_wr_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_data1=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_data[63:32]),UVM_HIGH)
			end

			else if(wb_trans_h.reg_addr==`TX2_ADDR) begin
				wb_trans_h.mon_data[95:64]=wb_trans_h.reg_wr_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_data2=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_data[95:64]),UVM_HIGH)
			end

			else if (wb_trans_h.reg_addr==`TX3_ADDR) begin
				wb_trans_h.mon_data[127:96]=wb_trans_h.reg_wr_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_data3=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_data[127:96]),UVM_HIGH)
			end
	
			if(wb_trans_h.reg_addr==`CTRL_STATUS_ADDR) begin
				cntrl_status_reg=wb_trans_h.reg_wr_data;
		//	`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h cntrl_status_reg=%h ",$time,wb_trans_h.reg_addr,cntrl_status_reg[31:0]),UVM_MEDIUM)
			end

		end

  		 else 
	 	 begin
			wb_trans_h.reg_addr <= wb_vif.wb_adr_i;
			wb_trans_h.reg_rd_data  = wb_vif.wb_dat_o;
			
			
			if(wb_trans_h.reg_addr==`RX0_ADDR) begin
				wb_trans_h.mon_rx_data[31:0]=wb_trans_h.reg_rd_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_rx_data0=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_rx_data[31:0]),UVM_HIGH)
				if(cntrl_status_reg[7:0]<=32) begin
					wb_analysis_port.write(wb_trans_h);
				end
			end


			else if(wb_trans_h.reg_addr==`RX1_ADDR) begin
				wb_trans_h.mon_rx_data[63:32]=wb_trans_h.reg_rd_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_rx_data1=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_rx_data[63:32]),UVM_HIGH)
				if(cntrl_status_reg[7:0] <=64 || cntrl_status_reg[7:0] > 32 ) begin
					wb_analysis_port.write(wb_trans_h);
				end
			end

			else if(wb_trans_h.reg_addr==`RX2_ADDR) begin
				wb_trans_h.mon_rx_data[95:64]=wb_trans_h.reg_rd_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_rx_data2=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_rx_data[95:64]),UVM_HIGH)
				if(cntrl_status_reg[7:0] <=96 || cntrl_status_reg[7:0] > 64 ) begin
					wb_analysis_port.write(wb_trans_h);
				end
			end

			else if (wb_trans_h.reg_addr==`RX3_ADDR) begin
				wb_trans_h.mon_rx_data[127:96]=wb_trans_h.reg_rd_data;
			`uvm_info(get_type_name(),$sformatf("*****[%0t] wb_trans_h.reg_addr=%h wb_trans_h.mon_rx_data3=%h ",$time,wb_trans_h.reg_addr,wb_trans_h.mon_rx_data[127:96]),UVM_HIGH)
				if(cntrl_status_reg[7:0] <=128 || cntrl_status_reg[7:0] > 96 ) begin
					wb_analysis_port.write(wb_trans_h);
				end
			end

		end
	//	`uvm_info(get_type_name(),$sformatf("[%0t]=============================================WB_MONITOR_from_dut ======================================= \n %s",$time,wb_trans_h.sprint()),UVM_MEDIUM)

	//scoreboard write method
		
	//	wb_analysis_port.write(wb_trans_h);
		end
	end

	`uvm_info("WB_MONITOR","WB_MONITOR_BEFORE_DROP_OBJECTION ", UVM_HIGH)
	phase.drop_objection(this);
 	`uvm_info("WB_MONITOR","WB_MONITOR_AFTER_DROP_OBJECTION ", UVM_HIGH)

 	  endtask : run_phase
endclass 



`include "reset_seq.sv"
`include "lsb_fst_data.sv"
`include "msb_fst_data_seq.sv"
`include "miso_data.sv"
